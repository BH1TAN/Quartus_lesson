module exp41(
			
			
			);
	
			